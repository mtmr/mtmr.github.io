network analysis example   
v1 1 0  
v2 3 0 dc 7    
r1 1 2 4      
r2 2 0 2
r3 2 3 1
.dc v1 28 28 1  
.print dc v(1,2) v(2,0) v(2,3)  
.end    


